`include "params.bsv"

typedef Bit#(INP_LEN) SysType;
typedef Bit#(INP_LEN * MAT_DIM) InpStreamType;
typedef Bit#(INP_LEN * MAT_DIM * MAT_DIM) OutStreamType;