`define STATE_DIM 6
`define INPUT_DIM 6
`define MEASUREMENT_DIM 2

`define INP_LEN 32
`define bits_int 16
`define bits_frac 16