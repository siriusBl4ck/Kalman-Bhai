`include "params.bsv"

typedef Bit#(INP_LEN) SysType;
typedef Bit#(INP_LEN * MAT_DIM) VecType;
typedef Bit#(INP_LEN * MAT_DIM * MAT_DIM) MatType;