`define INP_LEN 32
`define MAT_DIM 3
`define bits_int 16
`define bits_frac 16