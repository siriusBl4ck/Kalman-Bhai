package tb_mat_mult;

import mat_mult_systolic::*;

module tb_mat_mult(Empty);
    
endmodule

endpackage