`define INP_LEN 32
`define MAT_DIM 3